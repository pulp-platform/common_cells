
module cluster_level_shifter_in
(
    input  logic in_i,
    output logic out_o
);

assign out_o = in_i;

endmodule
