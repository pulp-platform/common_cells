
module pulp_level_shifter_out
  (
   input  logic in_i,
   output logic out_o
   );
   
   assign out_o = in_i;
   
endmodule
