/* Copyright (C) 2017 ETH Zurich, University of Bologna
 * All rights reserved.
 *
 * This code is under development and not yet released to the public.
 * Until it is released, the code is under the copyright of ETH Zurich and
 * the University of Bologna, and may contain confidential and/or unpublished 
 * work. Any reuse/redistribution is strictly forbidden without written
 * permission from ETH Zurich.
 *
 * Bug fixes and contributions will eventually be released under the
 * SolderPad open hardware license in the context of the PULP platform
 * (http://www.pulp-platform.org), under the copyright of ETH Zurich and the
 * University of Bologna.
 */

module pulp_clock_and2
(
    input  logic clk0_i,
    input  logic clk1_i,
    output logic clk_o
);

   C8T28SOI_LR_CNAND2X19_P0 ckand2
   (
      .Z(clk_o), 
      .A(clk0_i), 
      .B(clk1_i)
   );


endmodule
