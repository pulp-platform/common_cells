////////////////////////////////////////////////////////////////////////////////
// Company:        Multitherman Laboratory @ DEIS - University of Bologna     //
//                    Viale Risorgimento 2 40136                              //
//                    Bologna - fax 0512093785 -                              //
//                                                                            //
// Engineer:       Antonio Pullini - pullinia@iis.ee.ethz.ch                  //
//                                                                            //
// Additional contributions by:                                               //
//                                                                            //
//                                                                            //
//                                                                            //
// Create Date:    13/02/2013                                                 //
// Design Name:    ULPSoC                                                     //
// Module Name:    edge_propagator                                            //
// Project Name:   ULPSoC                                                     //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    edge_propagator                                            //
//                                                                            //
//                                                                            //
// Revision:                                                                  //
// Revision v0.1 - File Created                                               //
// Revision v0.2 - (19/03/2015)   clock_gating swapped in pulp_clock_gating   //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


module edge_propagator_tx
(
    input logic clk_i,
    input logic rstn_i,
    input logic valid_i,
    input logic ack_i,
    output logic valid_o
);

  reg [1:0] sync_a;
  
  reg  r_input_reg;
  wire s_input_reg_next;

  assign s_input_reg_next = valid_i | (r_input_reg & ~sync_a[0]);

  always @(negedge rstn_i or posedge clk_i)
  begin
    if (~rstn_i)
    begin
      r_input_reg <= 1'b0;
      sync_a      <= 2'b00;
    end
    else
    begin
      r_input_reg <= s_input_reg_next;
      sync_a      <= {ack_i,sync_a[1]};
    end
  end

  assign valid_o = r_input_reg;

endmodule








