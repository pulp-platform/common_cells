include/registers.svh